module dataPathMultiplier#(parameter N = 4)(
    output [N * 7 / 2 - 1:0] productDisp,
    input [N - 1:0] a,
    input [N - 1:0] b,
    input clk
);
    
endmodule
